library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is 
    Port ( address : in std_logic_vector(15 downto 0);
        write_data : in std_logic_vector(15 downto 0);
        MemWrite : in std_logic;
        read_data : out std_logic_vector(15 downto 0));
end memory;

architecture Behavioral of memory is
    type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);
    
    begin
        mem_process: process (address, write_data)
        
        variable data_mem : mem_array := (
        X"1201", -- LDR R0, =1
        X"1241", -- LDR R1, =1 
        X"1281", -- LDR R2, = 1
        X"0481", --ADI R2, R0, R1
        X"02C1", --ADD R3, R0, R1
        X"06D0", --INC R3, R2
        X"0881", --NOT R2, R0 
        X"0000", 
        X"0000", 
        X"0000", 
        X"0000",  
        X"0000",
        X"0000",  
        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000", X"0000",X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
        X"0000", X"0000");      
        
variable addr:integer;
begin -- the following type conversion function is in std_logic_arith
    addr:=conv_integer(address(8 downto 0));
    if MemWrite ='1' then
        data_mem(addr):= write_data;
    end if;
    --elsif MemRead='1' then
    read_data <= data_mem(addr) after 10 ns;
    --end if;
end process;
end Behavioral;